`timescale 1ns/10ps
module IIR_Real_testbench;
	parameter word_size_in = 64;
	parameter word_size_out = 2*word_size_in+2;
	parameter frac_bit = 52;

	reg [word_size_in-1:0] Data_in;
	reg clock, reset;
	wire [word_size_in-1:0] Data_out;

	IIR_Cheby1_Lowpass_Real DUT (
		.clock(clock),
		.reset(reset), 
		.Data_in(Data_in),
		.Data_out_r(Data_out)
	);

    initial 
    begin
        clock = 1'b0;
	    forever 
	    begin
			#10416 clock = ~clock;
			$display("At Time: %d  Filter Output=%d",$time,Data_out);
	    end  
    end

	initial
	begin
	  #0  reset=1;
		  Data_in=64'b0000000000000000000000000000000000000000000000000000000000000000;
	  #20832  reset=0;    
	  #20833  Data_in=64'b0000000000000010001101111100111011001011111000010101010000101110;
	  #20834  Data_in=64'b0000000000001000011001011100100110001000111010111001101011100010;
	  #20833  Data_in=64'b0000000000000100000110001001111110110011011111111110010111001011;
	  #20833  Data_in=64'b0000000000000001100010111010001101011000001110000101110000011100;
	  #20834  Data_in=64'b0000000000000000110000100001110101110010000000101001010100011101;
	  #20833  Data_in=64'b0000000000001001100110100010010000000111011100101100000101001101;
	  #20833  Data_in=64'b0000000000001000111100000101110011011110110100000100101100001000;
	  #20834  Data_in=64'b0000000000000110100000110111101101000100110010101000110110110011;
	  #20833  Data_in=64'b0000000000000110011000000100101011011100110001101001100010000001;
	  #20833  Data_in=64'b0000000000000110000110101101111100011011100100000001000100011111;
	  #20834  Data_in=64'b0000000000000110000101010100110110001001100111011000100101100000;
	  #20833  Data_in=64'b0000000000001001010110101001111010010111100100001100100010101001;
	  #20833  Data_in=64'b0000000000001001111110101001111100101010110101100000110101111000;
	  #20834  Data_in=64'b0000000000000001000000001011010101011010110100110100000101100000;
	  #20833  Data_in=64'b0000000000000000110101010101000100010110011111100110101110101101;
	  #20833  Data_in=64'b0000000000000100100111000000001110011011110100001110000101101100;
	  #20834  Data_in=64'b0000000000001000100101000110110110100100101101000111111001011110;
	  #20833  Data_in=64'b0000000000000010101010000010110011000001011000010000000011100000;
	  #20833  Data_in=64'b0000000000000000111001101001001100111101100100111100011110111010;
	  #20834  Data_in=64'b0000000000000001110100001010011001001001111100110001101000010101;
	  #20833  Data_in=64'b0000000000001000001010000100001111100000111001110110011001110010;
	  #20833  Data_in=64'b0000000000000011100010110100001010110101111110010000101111100010;
	  #20834  Data_in=64'b0000000000000010010000000111011011011111101000010011000110001011;
	  #20833  Data_in=64'b0000000000000000100011110011101111010100111110011010000100001111;
	  #20833  Data_in=64'b0000000000001001001010010001111100001010001100010000101110110010;
	  #20834  Data_in=64'b0000000000001000011111001100000000101011101111001110010001000101;
	  #20833  Data_in=64'b0000000000000110111010111001001010101001110100110001011010100010;
	  #20833  Data_in=64'b0000000000000110100101011100000100010101110001111101001000110100;
	  #20834  Data_in=64'b0000000000000101110001100001001111010010000011000000010101111011;
	  #20833  Data_in=64'b0000000000000101101000100110011011011001000100100011100000111101;
	  #20833  Data_in=64'b0000000000001001101110100011011010110100001111111001010011101101;
	  #20834  Data_in=64'b0000000000001010010010100001111011010010011010111010010100001110;
	  #20833  Data_in=64'b0000000000000001010010100011100011101000010111111000100010001010;
	  #20833  Data_in=64'b0000000000000000000111110000101111000010100110100101011110010110;
	  #20834  Data_in=64'b0000000000000101000101000010110011000100011100101011100001000100;
	  #20833  Data_in=64'b0000000000001000101101000000101111111010010101100110011011011110;
	  #20833  Data_in=64'b0000000000000011001000001010000110101010110011111001111100101010;
	  #20834  Data_in=64'b0000000000000001110010110111111100100110101101001111010111110001;
	  #20833  Data_in=64'b0000000000000001011100111011011001011100001011000001011101000101;
	  #20833  Data_in=64'b0000000000000111110111000010011010011000101011000111110010010111;
	  #20834  Data_in=64'b0000000000000010111101010100010111101111011100110001110100110100;
	  #20833  Data_in=64'b0000000000000010111100100100011000001011100000010110111010101111;
	  #20833  Data_in=64'b0000000000000000011010001011101011111001000000000000111101111100;
	  #20834  Data_in=64'b0000000000001000101010000010011111000001001001111111010010000111;
	  #20833  Data_in=64'b0000000000001000000000010010100110000111110111101110100111001100;
	  #20833  Data_in=64'b0000000000000111010011000100010001000111111101001101110101100011;
	  #20834  Data_in=64'b0000000000000110101110101101000011001100110000110011010010101101;
	  #20833  Data_in=64'b0000000000000101011000101010001010000110001001001100001110101010;
	  #20833  Data_in=64'b0000000000000101001011000010111011111011100101110010010000100100;
	  #20834  Data_in=64'b0000000000001010000011011110110001000101001010001111010111111101;
	  #20833  Data_in=64'b0000000000001010100010000101100000110001111110011000010010100110;
	  #20833  Data_in=64'b0000000000000001100111011011111101011001100011011101011000101101;
	  #20834  Data_in=64'b0000000000000000100101011001111010110110010100011100001111110100;
	  #20833  Data_in=64'b0000000000000101011111111111010000011010111010011011011011100111;
	  #20833  Data_in=64'b0000000000001000110001001010011000110111011001000001001000011110;
	  #20834  Data_in=64'b0000000000000011100111111111011001011110001001110100001011000010;
	  #20833  Data_in=64'b0000000000000010101011010010000000111111001010101010010010001101;
	  #20833  Data_in=64'b0000000000000001001000011110010001010100111100100000110100101000;
	  #20834  Data_in=64'b0000000000000111100000011110000010111010111001101101111101100001;
	  #20833  Data_in=64'b0000000000000010010110000001011100011110001110010010011001100111;
	  #20833  Data_in=64'b0000000000000011100111111001010011110010101011101111001000111101;
	  #20834  Data_in=64'b0000000000000000010011110010001101011010010101110101001011111100;
	  #20833  Data_in=64'b0000000000001000000101111111101001100001010000110010000100110010;
	  #20833  Data_in=64'b0000000000000111011111110000100011101111011000000110000010110110;
	  #20834  Data_in=64'b0000000000000111101001000101001000000100011001011001111001000011;
	  #20833  Data_in=64'b0000000000000110110011110010111100110100110011100111100011000101;
	  #20833  Data_in=64'b0000000000000100111100010110011001101110001010100110000110100010;
	  #20834  Data_in=64'b0000000000000100101101000001010001111111010010100110100110111101;
	  #20833  Data_in=64'b0000000000001010010101001001111100100011111000010010110011110010;
	  #20833  Data_in=64'b0000000000001010101101010010011111011110100111000110011100011011;
	  #20834  Data_in=64'b0000000000000001111110100100010000110110001001100110111110111000;
	  #20833  Data_in=64'b0000000000000001010001110010000111101011101110100110011001101001;
	  #20833  Data_in=64'b0000000000000101110111100100111111011010010111111101101001010001;
	  #20834  Data_in=64'b0000000000001000110001100110001111000111110110001100011110111101;
	  #20833  Data_in=64'b0000000000000100001001001101110111111010100100010111010101101000;
	  #20833  Data_in=64'b0000000000000011100010011101101010110001110110100010001111000101;
	  #20834  Data_in=64'b0000000000000000110110111111010110010100110011011101011011011100;
	  #20833  Data_in=64'b0000000000000111000110100000010110000000110000111011001100011110;
	  #20833  Data_in=64'b0000000000000001101101010011010100010001010100110111010111101010;
	  #20834  Data_in=64'b0000000000000100010001101111010011111011010001100001111111110001;
	  #20833  Data_in=64'b0000000000000000010000101101101000001001111001001000111011011100;
	  #20833  Data_in=64'b0000000000000111011110010111011000101000001100010101101111111011;
	  #20834  Data_in=64'b0000000000000110111101111101100110111001100001010000101101011000;
	  #20833  Data_in=64'b0000000000000111111100101001001001010101011010100100100010010100;
	  #20833  Data_in=64'b0000000000000110110100101011100001111000100010110111010000000110;
	  #20834  Data_in=64'b0000000000000100011100110101101001001010001111001100001110100010;
	  #20833  Data_in=64'b0000000000000100001110111000100100000101011011010000110011000000;
	  #20833  Data_in=64'b0000000000001010100011010100101011001111110110101010000011000110;
	  #20834  Data_in=64'b0000000000001010110100001001000111111011001111001000111000101100;
	  #20833  Data_in=64'b0000000000000010010111101010100111110111000001001011001001011101;
	  #20833  Data_in=64'b0000000000000001111100111111011011000001100011001100100010000010;
	  #20834  Data_in=64'b0000000000000110001011100101010111111010001001000111100000100111;
	  #20833  Data_in=64'b0000000000001000101110011001000101001111000000010000011010001001;
	  #20833  Data_in=64'b0000000000000100101011011111100100010011101010110011100001000000;
	  #20834  Data_in=64'b0000000000000100011000000001111000001101000101111111100111110110;
	  #20833  Data_in=64'b0000000000000000101000101000110110110111011010101000110010011010;
	  #20833  Data_in=64'b0000000000000110101001010100101100000111010100100111001011110000;
	  #20834  Data_in=64'b0000000000000001000011100010110000011101101101111111010111111100;
	  #20833  Data_in=64'b0000000000000100111001110000100001001111001100001110111000101101;
	  #20833  Data_in=64'b0000000000000000010001000001111110010011011010110010100110100111;
	  #20834  Data_in=64'b0000000000000110110011011001101101101001011101010011100101101110;
	  #20833  Data_in=64'b0000000000000110011011010001111011100111100110111100010011011001;
	  #20833  Data_in=64'b0000000000001000001101011111001101001010100001010111000100111010;
	  #20834  Data_in=64'b0000000000000110110001010111000000100110101000101100010111111110;
	  #20833  Data_in=64'b0000000000000011111010011001010111110010000100001111101010101011;
	  #20833  Data_in=64'b0000000000000011110000111111110110001000011101001000001000011010;
	  #20834  Data_in=64'b0000000000001010101101110000100100001001010000011110110010110001;
	  #20833  Data_in=64'b0000000000001010110110101100001000000101011111100100000100100101;
	  #20833  Data_in=64'b0000000000000010110010011011110011101100111010010001010101001111;
	  #20834  Data_in=64'b0000000000000010100110101001111100100101000101110001001010001010;
	  #20833  Data_in=64'b0000000000000110011011110011111001001111001000010100010100100001;
	  #20833  Data_in=64'b0000000000001000100111101001111111000011110000111000001011000100;
	  #20834  Data_in=64'b0000000000000101001110011101100100001100101101111000111101010110;
	  #20833  Data_in=64'b0000000000000101001011100110100011100011010101001001011011001010;
	  #20833  Data_in=64'b0000000000000000011101100010110100010101101011101101001110000001;
	  #20834  Data_in=64'b0000000000000110001001001000100010101101100010010011100001010100;
	  #20833  Data_in=64'b0000000000000000011001001001001001110010100111001011001001110100;
	  #20833  Data_in=64'b0000000000000101011111101000010100100101100001010010100111001101;
	  #20834  Data_in=64'b0000000000000000010100110000111100111111001000101001000011110001;
	  #20832  $stop;
	end

	
	initial 
	begin
		$dumpfile("IIR_dump.vcd");
		$dumpvars;
	end
endmodule
